module ALU #(parameter N=1) (
	input [N-1:0] a_i, b_i,
	input [3:0] ALUControl,
	output [N-1:0] y,
	output N_out, Z_out, C_out, V_out);
	

endmodule
