module testbenchFullAdder();

logic 
