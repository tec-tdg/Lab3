module testbenchFullAdder();





logic 
